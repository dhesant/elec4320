`include "define.v"

module alu(a, b, f, s);

 input [15:0] a, b;
 input [4:0] 	f;
 output [15:0] s;
 reg  [15:0] s;

//put your implementation here
//note: 'f' is the 5-bit opcode as in Table 2 in the manual.
//'a' and 'b' are the two operands

endmodule
